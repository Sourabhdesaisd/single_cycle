module ROL (

            input [31:0] in_1 ,
            input [31:0] in_2 ,

            output reg [31:0] out_rol

        ) ;

always@(*)
begin

    case(in_2[4:0])

        5'b00000 : out_rol = in_1;

        5'b00001 : out_rol = {in_1[30:0],in_1[31]};

        5'b00010 : out_rol = {in_1[29:0],in_1[31:30]};

        5'b00011 : out_rol = {in_1[28:0],in_1[31:29]};

        5'b00100 : out_rol = {in_1[27:0],in_1[31:28]};

        5'b00101 : out_rol = {in_1[26:0],in_1[31:27]};

        5'b00110 : out_rol = {in_1[25:0],in_1[31:26]};

        5'b00111 : out_rol = {in_1[24:0],in_1[31:25]};

        5'b01000 : out_rol = {in_1[23:0],in_1[31:24]};

        5'b01001 : out_rol = {in_1[22:0],in_1[31:23]};

        5'b01010 : out_rol = {in_1[21:0],in_1[31:22]};

        5'b01011 : out_rol = {in_1[20:0],in_1[31:21]};

        5'b01100 : out_rol = {in_1[19:0],in_1[31:20]};

        5'b01101 : out_rol = {in_1[18:0],in_1[31:19]};

        5'b01110 : out_rol = {in_1[17:0],in_1[31:18]};

        5'b01111 : out_rol = {in_1[16:0],in_1[31:17]};

        5'b10000 : out_rol = {in_1[15:0],in_1[31:16]};

        5'b10001 : out_rol = {in_1[14:0],in_1[31:15]};

        5'b10010 : out_rol = {in_1[13:0],in_1[31:14]};

        5'b10011 : out_rol = {in_1[12:0],in_1[31:13]};

        5'b10100 : out_rol = {in_1[11:0],in_1[31:12]};

        5'b10101 : out_rol = {in_1[10:0],in_1[31:11]};

        5'b10110 : out_rol = {in_1[9:0],in_1[31:10]};

        5'b10111 : out_rol = {in_1[8:0],in_1[31:9]};

        5'b11000 : out_rol = {in_1[7:0],in_1[31:8]};

        5'b11001 : out_rol = {in_1[6:0],in_1[31:7]};

        5'b11010 : out_rol = {in_1[5:0],in_1[31:6]};

        5'b11011 : out_rol = {in_1[4:0],in_1[31:5]};

        5'b11100 : out_rol = {in_1[3:0],in_1[31:4]};

        5'b11101 : out_rol = {in_1[2:0],in_1[31:3]};

        5'b11110 : out_rol = {in_1[1:0],in_1[31:2]};

        5'b11111 : out_rol = {in_1[0],in_1[31:1]};

    endcase

end

endmodule

